`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/20/2021 12:04:08 PM
// Design Name: 
// Module Name: serial_transmitter
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


//module serial_transmitter(
//    input clk,
//    output reg TX,
//    input [7:0] sending_buf,
//    output reg data_sent, //goes high when stop bit is sent
//    input [16:0] count_for_baud_rate,
//    input data_good
//);

//    reg [16:0] clock_count = 0;
//    reg currently_sending = 0;
//    reg [4:0] sent = 0;
//    reg enable = 0;
//    reg [7:0] sending = 0;
//    always@ (posedge clk) begin //sending in 8 bit chunks only for now
//        data_sent = 0;
//        clock_count <= clock_count + 1;
//        if(data_good) begin //reset state on aquisition of new data
//            sending <= sending_buf;
//            enable <= 1;
//            //sending_pos = 0;
//            //sent <= 0;
//            //currently_sending <= 0; 
//        end
//        if(clock_count == count_for_baud_rate) begin
//            clock_count <= 0;
//            if(currently_sending) begin //already sending byte
//                if(sent == 9) begin //need to finish byte with stop bit
//                    TX <= 1;
//                    sent <= 0;
//                    currently_sending <= 0;
//                    data_sent = 1;
//                end else begin //can continue with byte
//                    TX = sending[0];
//                    sending = sending >> 1;
//                    sent = sent + 1;
//                end
//            end else begin //starting new byte send with start bit
//                if(enable) begin//gates beginning of state machine behind enable
//                    TX <= 0;
//                    currently_sending <= 1;
//                    sent <= 1;
//                    enable <= 0;
//                end
//            end
//        end
//    end
//endmodule

module serial_transmitter #(parameter CLK_IN=0, parameter BAUD=0)( //no in built FIFO as of yet
    input clk,
    output reg TX,
    input wr_en, //is there new data on this clock edge
    output full,
    input [7:0] din,
    output [11:0] data_count//,
    //input [15:0] count_for_baud //max clock division of 2^16 -1
);
    parameter count_for_baud = CLK_IN / BAUD;
    
    import types::*;
    reg srst = 0; //I don't use reset at the moment
    reg rd_en = 0;

    wire empty;
    wire [7:0] dout;
    wire valid;
    uart_fifo fifo(
        .clk,
        .srst,
        .din,
        .wr_en,
        .rd_en,
        .dout,
        .full,
        .empty,
        .valid,
        .data_count
    );

    enum {WAITING='b00001, START_SENDING='b00010, DATA_SENDING='b00100, WAITING_AFTER_DATA='b01000, STOP_SENDING='b10000} current_state = WAITING;




    logic [15:0] clock_count = count_for_baud; //internal count to clock divide for proper baud rate
    logic [7:0] shift_reg = 0;

    logic [2:0] shift_pos = 0;



    always_ff @(posedge clk) begin
        case(current_state)
            WAITING: begin //send out a flag when it goes into waiting mode to see if this is duplicating characters
                TX <= 1;
                if(valid) begin
                    current_state <= START_SENDING;
                    shift_reg <= dout;
                    rd_en <= 1;
                end
            end
            START_SENDING: begin
                rd_en <= 0;
                TX <= 0;
                shift_pos <= 0;
                clock_count <= 0;
                current_state <= DATA_SENDING; //no delay needed here since DATA_SENDING starts instead of ends with a delay
            end
            DATA_SENDING: begin
                if(clock_count == count_for_baud) begin
                    clock_count <= 0;
                    TX <= shift_reg[shift_pos];
                    shift_pos <= shift_pos + 1;
                    if(shift_pos == 7)
                        current_state <= WAITING_AFTER_DATA;
                end else
                    clock_count <= clock_count + 1;
            end
            WAITING_AFTER_DATA: begin
                shift_reg <= 0;
                if(clock_count == count_for_baud) begin
                    clock_count <= 0;
                    current_state <= STOP_SENDING;
                end else
                    clock_count <= clock_count + 1;

            end
            STOP_SENDING: begin
                TX <= 1;
                if(clock_count == count_for_baud) begin
                    clock_count <= 0;
                    current_state <= valid ? START_SENDING : WAITING;
                    if(valid) begin
                        shift_reg <= dout;
                        rd_en <= 1;
                    end
                end else
                    clock_count <= clock_count + 1;
            end
            default: begin
                TX <= 1;
                current_state <= WAITING;
            end
        endcase
    end
    //    always_ff @(posedge clk) begin
    //        if((data_ready && !going) || (going && !data_ready)) begin //data_ready will interupt currently transmitting data for now
    //            if (clock_count == count_for_baud) begin
    //                clock_count <= '0;
    //                if(state_pos == 0) begin
    //                    going <= 1; //so that data_ready is only needed on the clock pulse the data is submitted
    //                    shift_reg <= data_ready ? data : shift_reg;
    //                    TX <= 0; //start bit
    //                    state_pos <= 1;
    //                    data_sent <= 0;
    //                    shift_pos <= 0;
    //                end else if (state_pos == 9) begin
    //                    TX <= 1; //stop bit
    //                    state_pos <= '0;
    //                    data_sent <= 1;
    //                    going <= 0;
    //                end else begin //only other state is sending data
    //                    TX <= shift_reg[shift_pos];
    //                    //shift_reg <= shift_reg >> 1;
    //                    state_pos <= state_pos + 1;
    //                    shift_pos <= shift_pos + 1;
    //                end

    //            end else begin
    //                clock_count <= clock_count + 1;
    //                data_sent <= '0;
    //            end
    //        end else begin
    //            if(data_ready)
    //                shift_reg <= data_ready;
    //            TX <= 1;
    //            data_sent <= 0;
    //            state_pos <= '0;
    //            clock_count <= count_for_baud; //make it go immediately
    //        end
    //    end
endmodule